module mult16bit_tb();
wire [31:0]t_p;
reg [15:0]t_a, t_b;

mult16bit my_multiplier_16(.a(t_a), .b(t_b), .p(t_p));
initial begin
$monitor("%d	%d	%d", t_a, t_b, t_p);

t_a=16'b10000001;
t_b=16'b11111111;
#100

t_a=16'b11001100;
t_b=16'b10101010;
#100

t_a=16'b10000111;
t_b=16'b11100011;
#100

t_a=16'b11000000;
t_b=16'b00000111;
#100

t_a=16'b1111111111111111;
t_b=16'b1111111111111111;
#100

t_a=16'b1111000011110000;
t_b=16'b1111010101010101;
#100

t_a=16'habcd;
t_b=16'b1001100110011001;
#100

t_a=16'b1101110111011101;
t_b=16'b1111111111111111;
#100

t_a=16'b0101000011110000;
t_b=16'b1001000011110000;
#100


t_a=16'b1000000000000000;
t_b=16'b1101110111011101;

end
endmodule
 
  
module booth16bit_tb();
wire [31:0]t_p;
reg [15:0]t_a, t_b;

booth16bit my_multiplier_16(.a(t_a), .b(t_b), .p(t_p));
initial begin
$monitor("a=%b	b=%b	p=%b", t_a, t_b, t_p);

t_a=16'sb1000000010011001;//-32615
t_b=16'sb1010101000000001;//22015
#100

t_a=-16'sd126;//-126
t_b=-16'sd1;//-1
#100

t_a=16'sb1000000011110101;//-32523
t_b=16'sb1010101001111000;//-21896
#100

t_a=16'sb0111111111111111;//-32767
t_b=16'sb0111111111111111;//-32767
#100

t_a=16'sb0101111010100110;//24230
t_b=16'sb0110110101011010;//27994
#100

t_a=16'sb1;//1
t_b=16'sb1;//1
#100

t_a=16'sh7a;//122
t_b=16'sb1000100100111001;//-30407
#100

t_a=16'sb0111011101111101;//30589
t_b=16'sb1010111110001111;//-20593
#100

t_a=16'sb1000001010100101;//-32091
t_b=-16'sb0111110000111001;//-31801
#100

t_a=-16'sb0101000001001100;//-20556
t_b=16'sb1000000010100101;//-32603

end
endmodule
 
  